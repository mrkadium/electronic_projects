��  CCircuit��  CSerializeHack           ��  CPart              ���  CLED�� 	 CTerminal  ����      	        �          
�  ����                            ����        ��      ��  CEarth
�  ���                            ��        ��      �� 	 CResistor��  CValue  `~��    0.16k   ������c@      �?k  
�  |���               �          
�  P�e�      	        �            d�|�        ��      ��  CAND
�  �p�q              @          
�  ����      	       @          
�  �x	y              @            �l��           ��    �� 	 CInverter
�  ����               �          
�  ����              @            �t��           ��    �
�  �@�A                          
�  �P�Q               �          
�  �H	I               �            �<�T            ��    ��  COR
�  XY               �          
�  hi              @          
�  4`Ia              @            T4l     %      ��    #�
�  �%�               �          
�  �%�               �          
�  <�Q�               �            $�<�     )      ��    �
�  �p�q              @          
�  ����               �          
�  �xy               �            �l��     -      ��    �
�  ����               �          
�  ����              @            ����     1      ��    �
�  ����               �          
�  ����      	       @          
�  ���               �            ����     4      ��    #�
�  %               �          
�   %!     
          �          
�  <Q               �            $<$     8      ��    �
�  ����              @          
�  ��	               �          
�  �                �            ���     <      ��    �
�  �8�9               �          
�  �8�9     	         @            �,�D     @      ��    �
�  �(�)                          
�  �8�9     	 	       @          
�  �01     
          �            �$�<     C      ��    ��  CBattery�  � � �     5V(          @      �? V 
�  � � !              @          
�  � � � �                              � � �     I    ��      ��  CSPST��  CToggle  P�p�      L   
�  @�U�              @          
�  l���               �            T�l�     O      ��    K�M�  `x��      Q   
�  Ppeq              @          
�  |p�q               �            dl|t     S      ��    �
�  � (� )                            � � 2    V    ��                    ���  CWire  ����      X�  H	Y       X�  h	y       X�  �P�Q      X�  ��       X�  x�       X�  ����      X�  H`Iq       X��� 
 CCrossOver  �$�,        ��9       X�   1      
 X�          X�  P�Q       X�  �8�9      X�  Hp�q      X�b�  ����        P���      X�  ��	      X�b�  �$�,      b�  �$�,        (�)      X�  @�A      X�b�  �l�t        �P��       X�  �  � q       X�b�  �l�t      b�  lt        � p�q      X�  � p� �       X�b�  ����      b�  ��        � ���      X�  � �A�      X�b�  ~d�l        �8��       X�  �8�9      X�b�  ����      b�  �$�,        ���9       X�  � h� �       X�  PhQq       X�b�  ����        ����       X�  ���q       X�b�  ~d�l        � hQi      X�b�  � $� ,        � �� i       X�b�  � $� ,        � ()      X�b�  ��      b�  lt        @)                     �                                 Y  Y      +   s       [  p       o   ! \ ! " " Z % Z % & [ & ' ' ` ) ^ ) * ] * + +  - h - . _ . / / ^ 1 � 1 2 2 5 4 i 4 5 2 5 6 6 ] 8 e 8 9 d 9 : : f < w < = k = > > e @ a @ A A D C l C D A D E E d I I r J   J O z O P P { S � S T T � V V �   " % &  p ! * 6 / ) � . ' h a m k g 9 E > 8 i : } @ ` - i � f 4 a = l c l � � C �   p t \ ~ I s s q s � v  r � w  w � v < � O { � } P { ~ ~ x ~ n  g � z � S � j _ � 1 T � | � � � � w � � � V � � y � u o l             �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 