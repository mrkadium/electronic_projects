��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  � "'    Enable (alta)      �  a�'    Enable (baja)      �  � �� �    	Selectora      �  � a� o    I0      �  � �� �    I1      �� 	 CGroupBox  � <��                           ���  CLogicIn�� 	 CLatchKey  (8'         �� 	 CTerminal  @$A9                            <D$        ����     ��  ��'        �  �$�9              @            ��$       ����     �� 	 CInverter�  �8�M       	       @          �  �d�y      	        �            �L�d          ��    ��  CAND�  @hUi              @          �  @xUy              @          �  lp�q              @            Tdl|           ��    ��  @�U�              @          �  @�U�     	 	        �          �  l���               �            T�l�     #      ��    ��   ��              @          �  ,�A�     	          �            �,�     '      ��    ��  � �� �     )   �  � �� �              @            � �� �     +   ����     ��  � a� o     ,   �  � h� i              @            � d� l     .   ����     ��  � �� �     /   �  � �� �               @            � �� �    1   ����     ��  COR�  ����              @          �  ����               �          �  ����              @            �|��     4      ��    ��  �x�y               �          �  ����      	       @          �  ���               �            �t��     8      ��    �� 	 CLogicOut�   ��      	        �            x$�     =      ��                  ���  CWire  � xAy      ?�  � ��      ?�  � hAi      ?��� 
 CCrossOver  � �� �        � �A�      ?�  � �� �       ?�D�  � �� �        � x� �       ?�  ����       ?�  �p��                     �                                        8  B    @   ! ! J # C # $ ( $ % % I ' A ' ( ( $ + + C . . B 1 F 1 4 J 4 5 I 5 6 6 9 8  8 9 6 9 : : = = : = G   F ' .  C H + # G 1 G E @ A 5 % ! 4             �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 