��  CCircuit��  CSerializeHack           ��  CPart              ���  CLogicIn�� 	 CLatchKey  ����     	   �� 	 CTerminal  ����              @            ����       ����     �� 	 CRailThru�  ����       d       @          �  ����      	       @            ����        ����    �
�  � � � �         �  � � � 	              @            � � � �        ����     ��  CAND�  8P9e      	          �          �  (P)e                �          �  0|1�               �            $d<|          ��    ��  H� ]�                �          �  H� ]�      	          �          �  t� ��                �            \� t�            ��    ��  CJK�  � �5                �          �  �8�9               �          �  �H�I              @          �  �X�Y               �          �  �\�q               �          �  �P�Q              @          �  �@�A               �            �4�\          ��   (   ��   5                �          �  �89               �          �  �HI              @          �  �XY               �          �  \q               �          �  $P9Q     
         @          �  $@9A     	          �            4$\     (    ��   (   ��  ` a5                �          �  @8U9              @          �  @HUI              @          �  @XUY              @          �  `\aq               �          �  tP�Q              @          �  t@�A               �            T4t\     0    ��   (                 ���  CWire  �� �A       8��� 
 CCrossOver  n�t�        pHq�       8�  p���      8�;�  n�t�        ���      8�  �@�A      8�  �@�A      8�  8� 9Q      	 8�  @� 9�      	 8�;�  >� D�         @� A�       	 8�;�  >� D�         �� I�       8�  8� A�      	 8�  @� I�      	 8�  xX�Y      8�;�  vD|L        x8yY       8�;�  vD|L        pH�I      8�  x8�9      8�  �� �9       8�  �� ��       8�  8� 9A      	 8�  �@�A      8�  �@�Y       8�;�  �T�\        �X�Y      8�;�  �T�\      ;�  ����        �H��       8�  �H�I      8�  (@)Q       8�  �@)A      8�;�  ����        `��      8�  p�       8�  ��1�      8�  �p��       8�  `pa�       8�  0HAI      8�;�  .T4\        0H1�       8�;�  .T4\        � XAY      8�  0���      8�  ��q�      8�  � 8� Y       8�  � 8A9      8�  � � 9       8�  �8�9      8�  �8�A                     �                               =       l  B   [    `  F   I    Q       ! P ! " M " # J # $ $ a % %   & & \ (   ( ) m ) * Z * + U + , , _ - -   . . R 0   0 1 k 1 2 c 2 3 f 3 4 4 b 5 5   6 6 A F S : ? M i :  > < ] a S n 6 9 C  D B D G C I F E 9  R D H  K # K N O J M L : " K ! Q O  P H . A T @ U U X T + W V W ^ Z i W * \  & [ ] Y b _ , > >  $ ` 4 ] d 2 d g c h f e j 3 d W h = k f l 1  j n ) m @            �%s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 