��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  � !� /    Set      �  � �� �    Reset      �  ����    Reset      �  ��    Set                    ��� 	 CLogicOut�� 	 CTerminal  ����              @            �x�          ��    ��  ��               �            �            ��    ��  CNAND�  �x�y               �          �  ����               �          �  ����              @            �t��           ��    ��  ��              @          �  � �!              @          �  ��               �            ��$           ��    ��  CSPDT��  CToggle   X@x         �  H%I      	       @          �  <PQQ               �          �  <@QA              @            $<<T            ��    ��  CBattery��  CValue  � /=    5V         @      �? V �  � HI              @          �  � H� I                            � <� T    '    ��      ��  `X�x     )   �  PHeI      	       @          �  |P�Q              @          �  |@�A     
          �            d<|T     +     ��    ��  `u              @            t�     /     ��    ��  CNOR�  ��	     
          �          �  ��     	          �          �  �              @            ��     2      ��    0��  �x�y              @          �  ����              @          �  ��     	          �            �t�     6      ��    ��  `�u�     	          �            tx��     :      ��    #�%�  /D=    5V         @      �? V �  <HQI              @          �  H%I               �            $<<T    =    ��      #�%�  d _� m    5V         @      �? V �  � x� y              @          �  X xm y                            l l� �    A    ��      ��  CSPST�  � �� �     D   �  � �� �              @          �  � �� �              @            � �� �     F     ��    C��  � @� `     H   �  � 8� 9              @          �  � 8� 9              @            � 4� <     J     ��    ��  ����              @            ����     M     ��    ��  �H�I               �            �@�P     O      ��    ��  `�u�               �          �  `�u�              @          �  ����              @            t���     Q      ��    ��  `@uA              @          �  `PuQ              @          �  �H�I               �            t<�T     U      ��    C��  ����     X   �  ����              @          �  ��	�              @            ����     Z     ��    C��  �@�`     \   �  �8�9              @          �  �89              @            �4�<     ^     ��    #�%�  |W�e    5V         @      �? V �  �p�q              @          �  pp�q                            �d�|    b    ��      ��  ����               �            ����     e      ��    0��  0�E�               �          �  0�E�              @          �  \�q�               �            D�\�     g      ��    0��  (8=9              @          �  (H=I               �          �  T@iA               �            <4TL     k      ��    ��  �@�A               �            �8�H     o      ��                  ���  CWire  ��      q�  ����      q�  �X��       q�  xx�y      q��� 
 CCrossOver  vT|\        xHyy       q�w�  vT|\        hX�Y      q�  xH�I      q�  ��I       q�  h iY       q�  h �!      q�  PPQ�       q�  P���      q�  PQA       q�  P�      q�  ����      q�  �P��       q�  �@�y       q�  ��	     
 q�  ��A      
 q�  0�      	 q�  �a�     	 q�w�  ,4        �01     	 q�  ��1      	 q�w�  ,4        A       q�  �@A      q�  a      q�  � 8� y       q�  � x� �       q�  � �� �      q�  � 8� 9      q�  � @aA      q�  � 8� A       q�  � �a�      q�  �H�I      q�  ����      q�  ����       q�  X�a�      q�w�  V�\�        XxY�       q�w�  V�\�        H���      q�  Xx�y      q�  �H�y       q�  HPaQ      q�  HPI�       q�   8)9      q�  �1�      q�  ����      q�  �p��       q�  �8�9      q�  �8�q       q�  h@�A      q�  0piq      q�w�  f\ld        h@iq       q�  (H)a       q�w�  f\ld        (`qa      q�  p���      q�  p`q�       q�  0p1�                     �                             s   r   u   �    t  �   ~    |   '   ! !  " " � ' '   (   ( + = + , , � - - � / � / 2 � 2 3 � 3 4 4 � 6 � 6 7 � 7 8 8 � : � : = = + >   > A A � B   B F � F G G � J � J K K � M � M O � O Q � Q R � R S S � U � U V � V W W � Z � Z [ [ � ^ � ^ _ _ � b b � c   c e � e g � g h � h i i � k � k l � l m m � o � o     y s v  v z { u y x } t v | r { ~ y }  ! �   � " �  � 7 , � � 6 � 2 � - � 8 � : � � � � 3 � � � � � � � 4 / � A � � � F � J � U K � G R W O S M � � � Q � � � � � � � � � � � � � V � � _ k [ h � Z b � � ^ � � m o � � � � � � l � � � � � � e � i � g             �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 